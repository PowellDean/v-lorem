module main

import lorem

fn main() {
    println(lorem.paragraphs(2))
}
